*SPICE LEVEL 2 PARAMETERS
 
.MODEL nenh nmos LEVEL=2 LD=0.181362U TOX=402.000000E-10
+ NSUB=6.567000E+15 VTO=0.805287 KP=4.757000E-05 GAMMA=0.5435
+ PHI=0.6 UO=553.83 UEXP=0.151038 UCRIT=48309.6
+ DELTA=0.823727 VMAX=50459.8 XJ=0.250000U LAMBDA=3.437039E-02
+ NFS=4.094390E+12 NEFF=1 NSS=1.000000E+12 TPG=1.000000
+ RSH=19.340000 CGDO=2.336825E-10 CGSO=2.336825E-10 CGBO=7.582249E-10
+ CJ=1.011600E-04 MJ=0.633000 CJSW=5.320000E-10 MJSW=0.266000 PB=0.800000
* Weff = Wdrawn - Delta_W
* The suggested Delta_W is 0.40 um
.MODEL penh pmos LEVEL=2 LD=0.250000U TOX=402.000000E-10
+ NSUB=6.786000E+15 VTO=-0.758994 KP=1.843000E-05 GAMMA=0.5525
+ PHI=0.6 UO=214.5 UEXP=0.253978 UCRIT=40136.1
+ DELTA=0.135535 VMAX=78961.6 XJ=0.050000U LAMBDA=4.876526E-02
+ NFS=4.352678E+11 NEFF=1.001 NSS=1.000000E+12 TPG=-1.000000
+ RSH=107.700000 CGDO=3.221216E-10 CGSO=3.221216E-10 CGBO=6.309201E-10
+ CJ=2.474000E-04 MJ=0.548900 CJSW=3.155000E-10 MJSW=0.327000 PB=0.800000
* Weff = Wdrawn - Delta_W
* The suggested Delta_W is -0.12 um
